*111
v1 1 0 10v
r1 1 0 20k
.control
run
print all
.endc
.end
* 课本 14章 例题 14.3.1 二极管电路

vi 1 0 PULSE(5v 0v 20us 0s 0s 10us 30us)

c1 1 2 CAP1 IC=0v
r1 2 0 10k
d1 3 2 DMOD
rl 3 0 10k

.model CAP1 C cap=50pf
.model DMOD D
.TRAN .1us 50us

.control
run
plot v(2) v(3)
.endc

.end

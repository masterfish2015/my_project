*tran 
v1 1 0 SIN(0 10v 50hz)

c1 1 2 20pf
r1 2 0 50Meg

.tran 1ms 20ms


.plot v(2)


.end
      

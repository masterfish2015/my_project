*exam 14.5.1
Vi  1 0 PWL(0 -1v 1s -1v 1.05s 1v 2s 1v 2.05s 3v 3s 3v)
Vcc 4 0 12V
Vtest_IB 2 99 0v

Rb  1 2 20k
Rc  4 3 3k

Q1  3 99 0 QMOD

.model QMOD NPN (BF=100)
.tran .01s 3s
.control
run
plot v(1) v(2) v(3)
plot -i(Vcc) vs i(Vtest_IB)
.endc
.end

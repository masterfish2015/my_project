* practice and think 14.3.7
v1 1 0 3v

*for test 
v_i_r2 2 99 0v

r1 1 2 1k
r2 99 0 1k

d1 2 0 DMOD

.model DMOD D

.op

.control
run
print all
.endc

.end
